module not_gate(a,y);
	input a;
	output y;
	not(y,a);
endmodule
