module or_gate(a,b,c);
	input a,b;
	output c;
	or(c,a,b);
endmodule
