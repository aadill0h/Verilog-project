module FCIMS_tb;

reg uprice0,uprice1,uprice2,uprice3,ncel0,ncel1,ncel2,ncel3,ct0,ct1,ct2,ct3,ctrl;
wire fprice0,fprice1,fprice2,fprice3,fprice4,fprice5,fprice6,fprice7,new_ct0,new_ct1,new_ct2,new_ct3;
FCIMS uut(ctrl,uprice0,uprice1,uprice2,uprice3,ncel0,ncel1,ncel2,ncel3,ct0,ct1,ct2,ct3,fprice0,fprice1,fprice2,fprice3,fprice4,fprice5,fprice6,fprice7,new_ct0,new_ct1,new_ct2,new_ct3);


initial begin
uprice0=0;uprice1=0;uprice2=0;uprice3=1;ncel0=1;ncel1=1;ncel2=0;ncel3=0;ct0=0;ct1=0;ct2=0;ct3=0;ctrl=0;
#10
uprice0=0;uprice1=0;uprice2=0;uprice3=1;ncel0=1;ncel1=1;ncel2=0;ncel3=0;ct0=1;ct1=1;ct2=0;ct3=0;ctrl=0;
#10
uprice0=0;uprice1=0;uprice2=0;uprice3=1;ncel0=0;ncel1=0;ncel2=1;ncel3=0;ct0=0;ct1=1;ct2=1;ct3=0;ctrl=1;
#10
$finish();
end
                
endmodule
